library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity demux is
    port (
        input:   in  std_logic;
        control: in  std_logic_vector(1 downto 0);
        output:  out std_logic_vector(3 downto 0)
    );
end demux;

architecture arch of demux is
    component and_gate is
        generic (
            N: natural := 3
        );

        port (
            input:  in  std_logic_vector(N - 1 downto 0);
            output: out std_logic
        );
    end component;

    component not_gate is
        port (
            input:  in  std_logic;
            output: out std_logic
        );
    end component;

    signal inv_control: std_logic_vector(1 downto 0);
begin
    -- for the inverse control
    u1: not_gate port map(control(0), inv_control(0));
    u2: not_gate port map(control(1), inv_control(1));

    u3: and_gate port map(inv_control                     & input, output(0));
    u4: and_gate port map(inv_control(1) &     control(0) & input, output(1));
    u5: and_gate port map(    control(1) & inv_control(0) & input, output(2));
    u6: and_gate port map(    control(1) &     control(0) & input, output(3));
end arch;

